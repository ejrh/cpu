module cpu(clk, do_reset);

    `include "parameters.v"
    
    input wire clk;
    input wire do_reset;

    wire do_fetch, do_regload, do_aluop, do_memload, do_memstore, do_regstore, do_next;
    
    wire [WORD_SIZE-1:0] pointer;
    wire [WORD_SIZE-1:0] pointer_adj;
    
    instr_pointer instr_pointer(pointer, pointer_adj, do_next, do_reset);

    wire [WORD_SIZE-1 : 0] instr;
    instr_fetch fetcher(instr, pointer, do_fetch);
    
    wire [NIB_SIZE-1 : 0] opcode, reg1, reg2, reg3;
    wire isaluop;
    wire [2 : 0] aluop;
    wire [BYTE_SIZE-1:0] bigval;
    wire [NIB_SIZE-1:0] smallval;
    instr_decode decoder(instr, opcode, isaluop, aluop, reg1, reg2, reg3, bigval, smallval);

    wire [WORD_SIZE-1 : 0] storeval, regval1, regval2;
    wire [NIB_SIZE-1 : 0] getnum1, getnum2, storenum;
    reg_stack stack(getnum1, getnum2, storenum, storeval, do_regload, do_regstore, regval1, regval2);
    
    wire get_sel;
    assign get_sel = (opcode == OP_STORE | opcode == OP_OUT
            | opcode == OP_BR | opcode == OP_LOADLO | opcode == OP_LOADHI);
    assign getnum1 = get_sel ? reg1 : reg2;
    assign getnum2 = get_sel ? reg2 : reg3;
    assign storenum = reg1;
    assign storeval = (opcode == OP_LOADLO) ? ((regval1 & 16'hFF00) | bigval)
            : (opcode == OP_LOADHI) ? ((regval1 & 16'h00FF) | (bigval << 8))
            : aluout;
    
    wire [WORD_SIZE-1 : 0] aluin1, aluin2;
    wire [WORD_SIZE-1 : 0] aluout;
    alu alu(aluop, aluin1, aluin2, do_aluop, aluout);
    
    assign aluin1 = regval1;
    assign aluin2 = regval2;

    reg [WORD_SIZE-1 : 0] reg1val, reg2val, reg3val;

    wire [0:WORD_SIZE-1] portaddr, portval;
    wire portget, portset;
    wire [0:WORD_SIZE-1] portout;
    ports ports1(portaddr, portval, portget, portset, portout);
    
    assign portaddr = regval2 + smallval;
    assign portval = regval1;
    assign portget = do_memload & (opcode == OP_IN);
    assign portset = do_memstore & (opcode == OP_OUT);
    
    control control(opcode, isaluop, clk, do_fetch, do_regload, do_aluop, do_memload, do_memstore, do_regstore, do_next);
    
    assign mux_adj = (opcode == OP_JMP) | (opcode == OP_BR & regval1 != 0);
    wire bigval_neg = bigval[BYTE_SIZE-1];
    assign pointer_adj = mux_adj ? (bigval_neg ? bigval - 256 : bigval) : 1;

endmodule
